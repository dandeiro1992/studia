LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY PC_1 IS PORT
(
A :IN STD_LOGIC_VECTOR(55 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
);
END PC_1;
--signal full_key:STD_LOGIC_VECTOR(63 DOWNTO 0):=A(55 downto 49) & '0' & A(48 downto 42) & '0' & A(41 downto 35) & '0' & A(34 downto 28) & '0' & A(27 downto 21) & '0' & A(20 downto 14) & '0' & A(13 downto 7) & '0' & A(6 downto 0) & '0';
ARCHITECTURE ARCH_PC_1 OF PC_1 IS
BEGIN
--Y(55)<=full_key(7);
--Y(54)<=full_key(15);
--Y(53)<=full_key(23);
--Y(52)<=full_key(31);
--Y(51)<=full_key(39);
--Y(50)<=full_key(47);
--Y(49)<=full_key(55);
--Y(48)<=full_key(63);
--Y(47)<=full_key(6);
--Y(46)<=full_key(14);
--Y(45)<=full_key(22);
--Y(44)<=full_key(30);
--Y(43)<=full_key(38);
--Y(42)<=full_key(46);
--Y(41)<=full_key(54);
--Y(40)<=full_key(62);
--Y(39)<=full_key(4);
--Y(38)<=full_key(13);
--Y(37)<=full_key(21);
--Y(36)<=full_key(29);
--Y(35)<=full_key(37);
--Y(34)<=full_key(45);
--Y(33)<=full_key(53);
--Y(32)<=full_key(61);
--Y(31)<=full_key(4);
--Y(30)<=full_key(12);
--Y(29)<=full_key(20);
--Y(28)<=full_key(28);
--Y(27)<=full_key(1);
--Y(26)<=full_key(9);
--Y(25)<=full_key(17);
--Y(24)<=full_key(25);
--Y(23)<=full_key(33);
--Y(22)<=full_key(41);
--Y(21)<=full_key(49);
--Y(20)<=full_key(57);
--Y(19)<=full_key(2);
--Y(18)<=full_key(10);
--Y(17)<=full_key(18);
--Y(16)<=full_key(26);
--Y(15)<=full_key(34);
--Y(14)<=full_key(42);
--Y(13)<=full_key(50);
--Y(12)<=full_key(58);
--Y(11)<=full_key(3);
--Y(10)<=full_key(11);
--Y(9)<=full_key(19);
--Y(8)<=full_key(27);
--Y(7)<=full_key(35);
--Y(6)<=full_key(43);
--Y(5)<=full_key(51);
--Y(4)<=full_key(59);
--Y(3)<=full_key(36);
--Y(2)<=full_key(44);
--Y(1)<=full_key(52);
--Y(0)<=full_key(60);

Y(55)<=A(6);
Y(54)<=A(13);
Y(53)<=A(20);
Y(52)<=A(27);
Y(51)<=A(34);
Y(50)<=A(41);
Y(49)<=A(48);
Y(48)<=A(55);
Y(47)<=A(5);
Y(46)<=A(12);
Y(45)<=A(19);
Y(44)<=A(26);
Y(43)<=A(33);
Y(42)<=A(40);
Y(41)<=A(47);
Y(40)<=A(54);
Y(39)<=A(4);
Y(38)<=A(11);
Y(37)<=A(18);
Y(36)<=A(25);
Y(35)<=A(32);
Y(34)<=A(39);
Y(33)<=A(46);
Y(32)<=A(53);
Y(31)<=A(3);
Y(30)<=A(10);
Y(29)<=A(17);
Y(28)<=A(24);
Y(27)<=A(0);
Y(26)<=A(7);
Y(25)<=A(14);
Y(24)<=A(21);
Y(23)<=A(28);
Y(22)<=A(35);
Y(21)<=A(42);
Y(20)<=A(49);
Y(19)<=A(1);
Y(18)<=A(8);
Y(17)<=A(15);
Y(16)<=A(22);
Y(15)<=A(29);
Y(14)<=A(36);
Y(13)<=A(43);
Y(12)<=A(50);
Y(11)<=A(2);
Y(10)<=A(9);
Y(9)<=A(16);
Y(8)<=A(23);
Y(7)<=A(30);
Y(6)<=A(37);
Y(5)<=A(44);
Y(4)<=A(51);
Y(3)<=A(31);
Y(2)<=A(38);
Y(1)<=A(45);
Y(0)<=A(52);
END ARCHITECTURE;