LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY PC_1 IS PORT
(
A :IN STD_LOGIC_VECTOR(55 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
);
END PC_1;
ARCHITECTURE ARCH_PC_1 OF PC_1 IS
signal full_key:STD_LOGIC_VECTOR(63 DOWNTO 0):=A(55 downto 49) & B"0" & A(48 downto 42) & B"0" & A(41 downto 35) & B"0" & A(34 downto 28) & B"0" & A(27 downto 21) & B"0" & A(20 downto 14) & B"0" & A(13 downto 7) & B"0" & A(6 downto 0) & B"0";
BEGIN
Y(55)<=full_key(7);
Y(54)<=full_key(15);
Y(53)<=full_key(23);
Y(52)<=full_key(31);
Y(51)<=full_key(39);
Y(50)<=full_key(47);
Y(49)<=full_key(55);
Y(48)<=full_key(63);
Y(47)<=full_key(6);
Y(46)<=full_key(14);
Y(45)<=full_key(22);
Y(44)<=full_key(30);
Y(43)<=full_key(38);
Y(42)<=full_key(46);
Y(41)<=full_key(54);
Y(40)<=full_key(62);
Y(39)<=full_key(5);
Y(38)<=full_key(13);
Y(37)<=full_key(21);
Y(36)<=full_key(29);
Y(35)<=full_key(37);
Y(34)<=full_key(45);
Y(33)<=full_key(53);
Y(32)<=full_key(61);
Y(31)<=full_key(4);
Y(30)<=full_key(12);
Y(29)<=full_key(20);
Y(28)<=full_key(28);
Y(27)<=full_key(1);
Y(26)<=full_key(9);
Y(25)<=full_key(17);
Y(24)<=full_key(25);
Y(23)<=full_key(33);
Y(22)<=full_key(41);
Y(21)<=full_key(49);
Y(20)<=full_key(57);
Y(19)<=full_key(2);
Y(18)<=full_key(10);
Y(17)<=full_key(18);
Y(16)<=full_key(26);
Y(15)<=full_key(34);
Y(14)<=full_key(42);
Y(13)<=full_key(50);
Y(12)<=full_key(58);
Y(11)<=full_key(3);
Y(10)<=full_key(11);
Y(9)<=full_key(19);
Y(8)<=full_key(27);
Y(7)<=full_key(35);
Y(6)<=full_key(43);
Y(5)<=full_key(51);
Y(4)<=full_key(59);
Y(3)<=full_key(36);
Y(2)<=full_key(44);
Y(1)<=full_key(52);
Y(0)<=full_key(60);
END ARCHITECTURE;