----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EXAMPLE IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE EXAMPLE_ARCH OF EXAMPLE IS
	COMPONENT schemat
	PORT
	(
		DATA_IN		:	 IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		CLK		:	 IN STD_LOGIC;
		DATA_OUT		:	 OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;
	TYPE MEMORY_BLOCK IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM : MEMORY_BLOCK;
	SIGNAL WEJSCIE :STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL WYJSCIE :STD_LOGIC_VECTOR(63 DOWNTO 0);
	
BEGIN
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (WR = '1') THEN
				MEM(conv_integer(ADDR)) <= DIN;
			ELSE
				WEJSCIE<=MEM(conv_integer(X"00000000")) & MEM(conv_integer(X"00000001"));
				MEM(conv_integer(X"00000002")) <= WYJSCIE(63 downto 32);
				MEM(conv_integer(X"00000003")) <= WYJSCIE(31 downto 0);
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(RD = '1') THEN
				DOUT <= MEM(conv_integer(ADDR));
			ELSE
				DOUT <= (others => 'Z');
			END IF;
		END IF;
	END PROCESS;
	
	--CEZAR1: entity work.Cezar port map(WEJSCIE(63 DOWNTO 0),WYJSCIE(63 DOWNTO 0));
	schem: schemat port map(DATA_IN=>WEJSCIE,CLK=>CLK,DATA_OUT=>WYJSCIE);
END ARCHITECTURE;