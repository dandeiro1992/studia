LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Przesuniecie IS PORT
(
DATA_IN :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
DATA_OUT :OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END Przesuniecie;
ARCHITECTURE ARCH_Przesuniecie OF Przesuniecie IS

BEGIN
DATA_OUT(7 downto 0)<=	X"44" WHEN DATA_IN(7 DOWNTO 0) =X"41"ELSE
								X"45" WHEN DATA_IN(7 DOWNTO 0) =X"42"ELSE
								X"46" WHEN DATA_IN(7 DOWNTO 0) =X"43"ELSE
								X"47" WHEN DATA_IN(7 DOWNTO 0) =X"44"ELSE
								X"48" WHEN DATA_IN(7 DOWNTO 0) =X"45"ELSE
								X"49" WHEN DATA_IN(7 DOWNTO 0) =X"46"ELSE
								X"4A" WHEN DATA_IN(7 DOWNTO 0) =X"47"ELSE
								X"4B" WHEN DATA_IN(7 DOWNTO 0) =X"48"ELSE
								X"4C" WHEN DATA_IN(7 DOWNTO 0) =X"49"ELSE
								X"4D" WHEN DATA_IN(7 DOWNTO 0) =X"4A"ELSE
								X"4E" WHEN DATA_IN(7 DOWNTO 0) =X"4B"ELSE
								X"4F" WHEN DATA_IN(7 DOWNTO 0) =X"4C"ELSE
								X"50" WHEN DATA_IN(7 DOWNTO 0) =X"4D"ELSE
								X"51" WHEN DATA_IN(7 DOWNTO 0) =X"4E"ELSE
								X"52" WHEN DATA_IN(7 DOWNTO 0) =X"4F"ELSE
								X"53" WHEN DATA_IN(7 DOWNTO 0) =X"50"ELSE
								X"54" WHEN DATA_IN(7 DOWNTO 0) =X"51"ELSE
								X"55" WHEN DATA_IN(7 DOWNTO 0) =X"52"ELSE
								X"56" WHEN DATA_IN(7 DOWNTO 0) =X"53"ELSE
								X"57" WHEN DATA_IN(7 DOWNTO 0) =X"54"ELSE
								X"58" WHEN DATA_IN(7 DOWNTO 0) =X"55"ELSE
								X"59" WHEN DATA_IN(7 DOWNTO 0) =X"56"ELSE
								X"5A" WHEN DATA_IN(7 DOWNTO 0) =X"57"ELSE
								X"41" WHEN DATA_IN(7 DOWNTO 0) =X"58"ELSE
								X"42" WHEN DATA_IN(7 DOWNTO 0) =X"59"ELSE
								X"43" WHEN DATA_IN(7 DOWNTO 0) =X"5A"ELSE
								(others=>'0');

END ARCHITECTURE;