LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.siphash_package.all;

ENTITY STER2 IS 
	PORT(	
	CLK	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	hash  :in  std_logic_vector(HASH_WIDTH-1 downto 0);
	
	DOUT     :out STD_LOGIC_VECTOR(31 downto 0)
	);
END ENTITY;

ARCHITECTURE rtl OF STER2 IS
	
	TYPE MEMORY_BLOCK IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM : MEMORY_BLOCK;

	
BEGIN
	

	PROCESS(CLK)
	BEGIN

	END PROCESS;
	
END ARCHITECTURE;