LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY iloczyn IS PORT
(
X :IN STD_LOGIC_VECTOR(1 DOWNTO 0);
Y :OUT STD_LOGIC
);
END ENTITY;

ARCHITECTURE arch_iloczyn OF iloczyn IS
BEGIN
Y <= (X(0) AND X(1));
END ARCHITECTURE;