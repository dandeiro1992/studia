----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EXAMPLE IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	RD   	:IN STD_LOGIC;
	WR		:IN STD_LOGIC;
	ADDR	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DIN	:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DOUT	:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE EXAMPLE_ARCH OF EXAMPLE IS
	
	--TYPE MEMORY_BLOCK IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	--SIGNAL MEM : MEMORY_BLOCK;
	
	SIGNAL PLAINTEXT :STD_LOGIC_VECTOR(63 DOWNTO 0):=X"0000000000000000";
	SIGNAL CIPHERTEXT :STD_LOGIC_VECTOR(63 DOWNTO 0):=X"0000000000000000";
	--SIGNAL BEGIN_NUMBER :STD_LOGIC_VECTOR(63 DOWNTO 0);
	--SIGNAL KEY		: STD_LOGIC_VECTOR(55 DOWNTO 0);
	SIGNAL STATE: STD_LOGIC:='0';
	SIGNAL END_FLAG:STD_LOGIC:='0';
	SIGNAL COMPARE_FLAG:STD_LOGIC:='0';
	SIGNAL COMPARE:STD_LOGIC:='0';
	SIGNAL END_NUMBER :STD_LOGIC_VECTOR(63 DOWNTO 0):=X"0000000000000000";
	SIGNAL COUNTER :STD_LOGIC_VECTOR(63 DOWNTO 0):=X"0000000000000000";
	SIGNAL RESULT		: STD_LOGIC_VECTOR(63 DOWNTO 0):=X"0000000000000000";
	SIGNAL FOUND_KEY:STD_LOGIC_VECTOR(55 DOWNTO 0):=X"00000000000000";
	
BEGIN
	PROCESS (CLK)
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			IF((ADDR(3 DOWNTO 0)=b"0000") AND (WR='1')) THEN
				PLAINTEXT(63 DOWNTO 32)<= DIN;
			END IF;
			IF((ADDR(3 DOWNTO 0)=b"0001") AND (WR='1')) THEN
				PLAINTEXT(31 DOWNTO 0)<= DIN;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (CLK)
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			IF((ADDR(3 DOWNTO 0)=b"0010") AND (WR='1')) THEN
				CIPHERTEXT(63 DOWNTO 32)<= DIN;
			END IF;
			IF((ADDR(3 DOWNTO 0)=b"0011") AND (WR='1')) THEN
				CIPHERTEXT(31 DOWNTO 0)<= DIN;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (CLK)
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			IF((ADDR(3 DOWNTO 0)=b"0100") AND (WR='1')) THEN
				COUNTER(63 DOWNTO 32)<= DIN;
			ELSIF((ADDR(3 DOWNTO 0)=b"0101") AND (WR='1')) THEN
				COUNTER(31 DOWNTO 0)<= DIN;
			ELSIF(STATE='1') THEN
				COUNTER(63 DOWNTO 8)<= std_logic_vector(unsigned(COUNTER(63 DOWNTO 8))+1);
			ELSE
				COUNTER<=COUNTER;	
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (CLK)
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			IF((ADDR(3 DOWNTO 0)=b"0110") AND (WR='1')) THEN
				END_NUMBER(63 DOWNTO 32)<= DIN;
			END IF;
			IF((ADDR(3 DOWNTO 0)=b"0111") AND (WR='1')) THEN
				END_NUMBER(31 DOWNTO 0)<= DIN;
			END IF;
		END IF;
	END PROCESS;

	PROCESS (CLK)
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			CASE STATE IS
				WHEN '0'=>
					IF(END_NUMBER(5)='1' AND COMPARE='0') THEN
						STATE<='1';
					ELSE
						STATE<='0';
					END IF;
				WHEN '1'=>
					IF(END_FLAG='1' OR END_NUMBER(4)='1' OR COMPARE='1') THEN
						STATE<='0';	
						--END_NUMBER(5)<='0';
					ELSE
						STATE<='1';
						--FOUND_KEY<=COUNTER(63 DOWNTO 8);
					END IF;
				when others => STATE<='0';
			END CASE;
		END IF;
	END PROCESS;
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(ADDR(3 DOWNTO 0)=b"1000" AND RD = '1') THEN
				DOUT <= FOUND_KEY(55 DOWNTO 28) & b"0000";
			ELSIF (ADDR(3 DOWNTO 0)=b"1000" AND RD = '1') THEN
				DOUT <= FOUND_KEY(27 DOWNTO 0) & b"0000";
			ELSE
				DOUT <= (others => 'Z');
			END IF;
		END IF;
	END PROCESS;
	
	
	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			if(COMPARE_FLAG='1') THEN
				COMPARE<='1';
			END IF;
		END IF;
	END PROCESS;
	
	
	--KEY <=CIPHERTEXT(63 DOWNTO 8);
	DES: entity work.des port map(PLAINTEXT,COUNTER(63 DOWNTO 8),RESULT);
	--done: entity work.DONE port map(CLK,BEGIN_NUMBER,CIPHERTEXT,END_NUMBER,PLAINTEXT,START,RESULT);
	
	END_FLAG<= '1' WHEN COUNTER=END_NUMBER(63 DOWNTO 8) ELSE '0';
	COMPARE_FLAG<='1'  WHEN (CIPHERTEXT=RESULT ) ELSE '0';
	FOUND_KEY<=COUNTER(63 DOWNTO 8);
END ARCHITECTURE;


