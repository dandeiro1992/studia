LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY COUNTER IS PORT(
BEGIN_NUMBER :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
END_NUMBER :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
COMPARISON_RESULT :IN STD_LOGIC;
CLK :IN STD_LOGIC;
NUMBER_OUT : OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
);
END COUNTER;

ARCHITECTURE ARCH_COUNTER OF COUNTER IS

SIGNAL START_NUMBER :STD_LOGIC_VECTOR (63 DOWNTO 0);
SIGNAL FINISH_NUMBER :STD_LOGIC_VECTOR (63 DOWNTO 0);
SIGNAL COUNTER :STD_LOGIC_VECTOR (55 DOWNTO 0);
SIGNAL FLAG: STD_LOGIC;

BEGIN

PROCESS(CLK)
	BEGIN
		IF(CLK'EVENT AND CLK='1') THEN
			IF(FINISH_NUMBER(2)='1') THEN
				COUNTER<=START_NUMBER(63 DOWNTO 8);
			ELSIF (FINISH_NUMBER(4)='1') THEN
				NUMBER_OUT<=COUNTER;
			ELSIF (FINISH_NUMBER(5)='1') THEN
				COUNTER<=std_logic_vector(unsigned(COUNTER)+1);
				NUMBER_OUT<=COUNTER;
			ELSE
				NUMBER_OUT<=COUNTER;
			END IF;
		END IF;
END PROCESS;

START_NUMBER <= BEGIN_NUMBER(63 DOWNTO 0);
FINISH_NUMBER(63 DOWNTO 5) <= END_NUMBER(63 DOWNTO 5);
FINISH_NUMBER(3 DOWNTO 0) <= END_NUMBER(3 DOWNTO 0);
FLAG<='1' WHEN COUNTER=END_NUMBER(63 DOWNTO 8) ELSE '0';
FINISH_NUMBER(4) <=COMPARISON_RESULT OR FLAG;
END ARCHITECTURE;
