LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY key_xor IS PORT
(
A :IN STD_LOGIC_VECTOR(47 DOWNTO 0);--nowo powstały podciag bitów
key :IN STD_LOGIC_VECTOR(47 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
);
END key_xor;

ARCHITECTURE ARCH_key_xor OF key_xor IS

BEGIN
Y<=A xor key;
END ARCHITECTURE;