LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Comparator IS PORT
(
CLK	:IN STD_LOGIC;
DATA_IN_1 :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
DATA_IN_2 :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
DATA_IN_3 :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
DATA_OUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END Comparator;
ARCHITECTURE ARCH_Comparator OF Comparator IS

BEGIN

	PROCESS(CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF(DATA_IN_1=DATA_IN_2) THEN
				DATA_OUT<=DATA_IN_1;
			ELSIF (DATA_IN_1=DATA_IN_3) THEN
				DATA_OUT<=DATA_IN_1;
			ELSIF (DATA_IN_2=DATA_IN_3) THEN
				DATA_OUT<=DATA_IN_2;
			ELSE 
				DATA_OUT<=(OTHERS=>'0');
			END IF;
		END IF;
	END PROCESS;
	
END ARCHITECTURE;