LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY work;

ENTITY DONE IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		BEGIN_NUMBER :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		CIPHERTEXT :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		END_NUMBER :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		PLAINTEXT :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		RESULT :  OUT  STD_LOGIC_VECTOR(55 DOWNTO 0)
	);
END DONE;

ARCHITECTURE bdf_type OF DONE IS 

COMPONENT des
	PORT(DATA_IN : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 KEY : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

COMPONENT counter
	PORT(COMPARISON_RESULT : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 BEGIN_NUMBER : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 END_NUMBER : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 NUMBER_OUT : OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
	);
END COMPONENT;

COMPONENT comparator
	PORT(CIPHERTEXT : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 DES_OUT : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		 KEY : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
		 COMPARISON_RESULT : OUT STD_LOGIC;
		 KEY_OUT : OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(55 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(63 DOWNTO 0);


BEGIN 

b2v_inst1 : counter
PORT MAP(COMPARISON_RESULT => SYNTHESIZED_WIRE_1,
		 CLK => CLK,
		 BEGIN_NUMBER => BEGIN_NUMBER,
		 END_NUMBER => END_NUMBER,
		 NUMBER_OUT => SYNTHESIZED_WIRE_4);
		 
b2v_inst : des
PORT MAP(DATA_IN => PLAINTEXT,
		 KEY => SYNTHESIZED_WIRE_4,
		 DATA_OUT => SYNTHESIZED_WIRE_2);

b2v_inst2 : comparator
PORT MAP(CIPHERTEXT => CIPHERTEXT,
		 DES_OUT => SYNTHESIZED_WIRE_2,
		 KEY => SYNTHESIZED_WIRE_4,
		 COMPARISON_RESULT => SYNTHESIZED_WIRE_1,
		 KEY_OUT => RESULT);


END bdf_type;